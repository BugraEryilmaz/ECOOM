`define LOG(x) $display x