// `define LOG(x) $display x
`define LOG(x) noAction
// `define debug 0