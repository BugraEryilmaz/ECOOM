`define LOG(x) $display x
`define debug 1